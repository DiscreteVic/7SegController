
module 7SegController(input [3:0]dig, input dot, output [7:0]leds);



	


endmodule
